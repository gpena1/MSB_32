///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: ALU_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Inputs: A (32-bit)
//         B (32-bit)
//         H (5-bit)
//         alu_op (7-bits: Shift, Ainvert, Binvert, CarryIn, Op2, Op1, Op0)
reg[31:0] A;
reg[31:0] B;
reg[4:0] H;
reg[6:0] alu_op;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Outputs: Result (32-bit)
//          Zero (1-bit)
//          Overflow (1-bit)
wire[31:0] Result;
wire zero;
wire overflow;
///////////////////////////////////////////////////////////////////////////////////

ALU_32 myALU(.A(A), .alu_op(alu_op), .B(B), .H(H), .Zero(zero), .Overflow(overflow), .Result(Result));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 & 21 = 5
$display("Testing: 45 & 21 = 5");
A=45; alu_op=7'b0000000; B=21;   #10; 
verifyEqual32(Result, A&B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 | 21 = 61
$display("Testing: 45 | 21 = 61");
A=45; alu_op=7'b0000001; B=21;   #10; 
verifyEqual32(Result, A|B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 + 21 = 66
$display("Testing: 45 + 21 = 66");
A=45; alu_op=7'b0000010; B=21;   #10; 
verifyEqual32(Result, A+B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 - 21 = 24
$display("Testing: 45 - 21 = 24");
A=45; alu_op=7'b0011010; B=21;   #10; 
verifyEqual32(Result, A-B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 < 21 = 0
$display("Testing: 45 < 21 = 0");
A=45; alu_op=7'b0011011; B=21;   #10; 
verifyEqual32(Result, A<B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 21 < 45 = 1
$display("Testing: 21 < 45 = 0");
A=21; alu_op=7'b0011011; B=45;   #10; 
verifyEqual32(Result, A<B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 NOR 21 = 2
$display("Testing: 45 NOR 21 = 2");
A=45; alu_op=7'b0110000; B=21;   #10; 
verifyEqual32(Result, ~(A|B));
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 NAND 21 = 58
$display("Testing: 45 NAND 21 = 58");
A=45; alu_op=7'b0110001; B=21;   #10; 
verifyEqual32(Result, ~(A&B));
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 == 21 = 0
A=45; alu_op=7'b0011010; B=21;   #10; 
$display("Testing if 45 == 21: 0");
verifyEqual(zero, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 == 45 = 1
A=45; alu_op=7'b0011010; B=45;   #10; 
$display("Testing if 45 == 45: 1");
verifyEqual(zero, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)+1 overflows
$display("Testing if (2^31-1)+1 overflows: 1");
A = 2147483647; B = 1; alu_op=7'b0000010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)+(-1) overflows
$display("Testing if (-2^31)+(-1) overflows: 1");
A = -2147483648; B = -1; alu_op=7'b0000010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)-1 overflows
$display("Testing if (-2^31)-1 overflows: 1");
A = -2147483648; B = 1; alu_op=7'b0011010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)-(-1) overflows
$display("Testing if (2^31-1)-(-1) overflows: 1");
A = 2147483647; B = -1; alu_op=7'b0011010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)<(-1) overflows (it will, < uses -)
$display("Testing if (2^31-1)<(-1) overflows: 1");
A = 2147483647; B = -1; alu_op=7'b0011011; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)<(1) overflows (it will, < uses -)
$display("Testing if (-2^31)<(1) overflows: 1");
A = -2147483648; B = 1; alu_op=7'b0011011; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 << 2 = 180
$display("Testing: 45 << 2 = 180");
B=45; H=2; alu_op=7'b1000000;   #10; 
verifyEqual32(Result, B*4);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 * 2 = 90
$display("Testing: 45 * 2 = 90");
A=45; B=2; alu_op=7'b0000100;   #10; 
verifyEqual32(Result, A*B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(0) = 0
$display("Testing: log2(0) = 0");
A=0; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(1) = 0
$display("Testing: log2(1) = 0");
A=1; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(2) = 1
$display("Testing: log2(2) = 1");
A=2; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(3) = 1
$display("Testing: log2(3) = 1");
A=3; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(4) = 2
$display("Testing: log2(4) = 2");
A=4; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 2);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(7) = 2
$display("Testing: log2(7) = 2");
A=7; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 2);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(8) = 3
$display("Testing: log2(8) = 3");
A=8; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 3);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(16) = 4
$display("Testing: log2(16) = 4");
A=16; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 4);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(31) = 4
$display("Testing: log2(31) = 4");
A=31; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 4);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(32) = 5
$display("Testing: log2(32) = 5");
A=32; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 5);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(1023) = 9
$display("Testing: log2(1023) = 9");
A=1023; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 9);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(1024) = 10
$display("Testing: log2(1024) = 10");
A=1024; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 10);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(2^31-1) = 30
$display("Testing: log2(2^31-1) = 30");
A=2147483647; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 30);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(2^31) = 31
$display("Testing: log2(2^31) = 31");
A=32'h80000000; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 31);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: log2(2^32-1) = 31
$display("Testing: log2(2^32-1) = 31");
A=32'hFFFFFFFF; alu_op=7'b0000011; B=0;   #10;
verifyEqual32(Result, 31);
////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
