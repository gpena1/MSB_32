///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: ALU_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Inputs: A (32-bit)
//         B (32-bit)
//         alu_op (5-bits: Ainvert, Binvert, CarryIn, Op1, Op0)
reg[31:0] A;
reg[31:0] B;
reg[4:0] alu_op;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Outputs: S (32-bit)
//          eq (1-bit)
//          overflow (1-bit)
wire[31:0] S;
wire zero;
wire overflow;
///////////////////////////////////////////////////////////////////////////////////

ALU_32 myALU(.A(A), .alu_op(alu_op), .B(B), .Overflow(overflow), .Zero(zero), .Result(S));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 & 21 = 5
$display("Testing: 45 & 21 = 5");
A=45; alu_op=5'b00000; B=21;   #10; 
verifyEqual32(S, A&B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 | 21 = 61
$display("Testing: 45 | 21 = 61");
A=45; alu_op=5'b00001; B=21;   #10; 
verifyEqual32(S, A|B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 + 21 = 66
$display("Testing: 45 + 21 = 66");
A=45; alu_op=5'b00010; B=21;   #10; 
verifyEqual32(S, A+B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 - 21 = 24
$display("Testing: 45 - 21 = 24");
A=45; alu_op=5'b01110; B=21;   #10; 
verifyEqual32(S, A-B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 < 21 = 0
$display("Testing: 45 < 21 = 0");
A=45; alu_op=5'b01111; B=21;   #10; 
verifyEqual32(S, A<B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 21 < 45 = 1
$display("Testing: 21 < 45 = 0");
A=21; alu_op=5'b01111; B=45;   #10; 
verifyEqual32(S, A<B);
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 NOR 21 = 2
$display("Testing: 45 NOR 21 = 2");
A=45; alu_op=5'b11000; B=21;   #10; 
verifyEqual32(S, ~(A|B));
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 NAND 21 = 58
$display("Testing: 45 NAND 21 = 58");
A=45; alu_op=5'b11001; B=21;   #10; 
verifyEqual32(S, ~(A&B));
$display("  Ensuring no overflow");
verifyEqual(overflow, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 == 21 = 0
A=45; alu_op=5'b01110; B=21;   #10; 
$display("Testing if 45 == 21: 0");
verifyEqual(zero, 0);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: 45 == 45 = 1
A=45; alu_op=5'b01110; B=45;   #10; 
$display("Testing if 45 == 45: 1");
verifyEqual(zero, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)+1 overflows
$display("Testing if (2^31-1)+1 overflows: 1");
A = 2147483647; B = 1; alu_op=5'b00010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)+(-1) overflows
$display("Testing if (-2^31)+(-1) overflows: 1");
A = -2147483648; B = -1; alu_op=5'b00010; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)-1 overflows
$display("Testing if (-2^31)-1 overflows: 1");
A = -2147483648; B = 1; alu_op=5'b01110; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)-(-1) overflows
$display("Testing if (2^31-1)-(-1) overflows: 1");
A = 2147483647; B = -1; alu_op=5'b01110; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (2^31-1)<(-1) overflows (it will, < uses -)
$display("Testing if (2^31-1)<(-1) overflows: 1");
A = 2147483647; B = -1; alu_op=5'b01111; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: (-2^31)<(1) overflows (it will, < uses -)
$display("Testing if (-2^31)<(1) overflows: 1");
A = -2147483648; B = 1; alu_op=5'b01111; #10;
verifyEqual(overflow, 1);
////////////////////////////////////////////////////////////////////////////////////////


$display("All tests passed.");
end

endmodule